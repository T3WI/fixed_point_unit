`timescale 1ns/1ps

module my_fpu_sim;
    
endmodule