package fpu_package;
    typedef enum {LOGIC_SHIFT, ARITH_SHIFT, CIRC_SHIFT, LZD, BARREL, REV, ADD, SUB, MUL, DIV,
    MAC} sel_modes;
endpackage